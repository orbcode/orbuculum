module time_stamp
(
  output wire [31:0]  time_dout
);
  assign time_dout  = 32'h5737ADFF;
endmodule
